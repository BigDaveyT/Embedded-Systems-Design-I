
module nios_system (
	clk_clk,
	leds_export_export,
	pushbuttons_export_export,
	reset_reset_n);	

	input		clk_clk;
	output	[7:0]	leds_export_export;
	input	[3:0]	pushbuttons_export_export;
	input		reset_reset_n;
endmodule
